/*
*
* Copyright (c) 2011 fpgaminer@bitcoin-mining.com
*
*
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published by
* the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
*
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <http://www.gnu.org/licenses/>.
* 
*/


`timescale 1ns/1ps

module e0 (x, y);

  input [31:0] x;
  output [31:0] y;

  assign y = {x[1:0],x[31:2]} ^ {x[12:0],x[31:13]} ^ {x[21:0],x[31:22]};

endmodule


module e1 (x, y);

  input [31:0] x;
  output [31:0] y;

  assign y = {x[5:0],x[31:6]} ^ {x[10:0],x[31:11]} ^ {x[24:0],x[31:25]};

endmodule


module ch (x, y, z, o);

  input [31:0] x, y, z;
  output [31:0] o;

  assign o = z ^ (x & (y ^ z));

endmodule


module maj (x, y, z, o);

  input [31:0] x, y, z;
  output [31:0] o;

  assign o = (x & y) | (z & (x | y));

endmodule


module s0 (x, y);

  input [31:0] x;
  output [31:0] y;

  assign y[31:29] = x[6:4] ^ x[17:15];
  assign y[28:0] = {x[3:0], x[31:7]} ^ {x[14:0],x[31:18]} ^ x[31:3];

endmodule


module s1 (x, y);

  input [31:0] x;
  output [31:0] y;

  assign y[31:22] = x[16:7] ^ x[18:9];
  assign y[21:0] = {x[6:0],x[31:17]} ^ {x[8:0],x[31:19]} ^ x[31:10];

endmodule


